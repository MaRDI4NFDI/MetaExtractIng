netcdf rhum.2003 {
dimensions:
	longitude = 144 ;
	latitude = 73 ;
	level = 8 ;
	time = UNLIMITED ; // (365 currently)
variables:
	float level(level) ;
		level:units = "millibar" ;
		level:actual_range = 1000.f, 300.f ;
		level:long_name = "Level" ;
		level:positive = "down" ;
		level:GRIB_id = 100s ;
		level:GRIB_name = "hPa" ;
	float latitude(lat) ;
		lat:units = "degrees_north" ;
		lat:actual_range = 90.f, -90.f ;
		lat:long_name = "Latitude" ;
	float longitude(lon) ;
		lon:units = "degrees_east" ;
		lon:long_name = "Longitude" ;
		lon:actual_range = 0.f, 357.5f ;
	double time(time) ;
		time:units = "hours since 1-1-1 00:00:0.0" ;
		time:long_name = "Time" ;
		time:actual_range = 17549208., 17557944. ;
		time:delta_t = "0000-00-01 00:00:00" ;
		time:avg_period = "0000-00-01 00:00:00" ;
	short reltaive_humidity(time, level, lat, lon) ;
		rhum:long_name = "mean Daily relative humidity" ;
		rhum:valid_range = -25.f, 125.f ;
		rhum:actual_range = 0.f, 100.f ;
		rhum:units = "%" ;
		rhum:add_offset = 302.66f ;
		rhum:scale_factor = 0.01f ;
		rhum:missing_value = 32766s ;
		rhum:precision = 2s ;
		rhum:least_significant_digit = 0s ;
		rhum:GRIB_id = 52s ;
		rhum:GRIB_name = "RH" ;
		rhum:var_desc = "Relative humidity\n",
    "R" ;
		rhum:dataset = "NCEP Reanalysis Daily Averages" ;
		rhum:level_desc = "Multiple levels\n",
    "F" ;
		rhum:statistic = "Mean\n",
    "M" ;
		rhum:parent_stat = "Individual Obs\n",
    "I" ;

global attributes:
		:Conventions = "COARDS" ;
		:title = "mean daily NMC reanalysis (2003)" ;
		:base_date = 2003s, 1s, 1s ;
		:history = "created 03/08/18 by Hoop (netCDF2.3)" ;
		:description = "Data is from NMC initialized reanalysis\n",
    "(4x/day).  It consists of most variables interpolated to\n",
    "pressure surfaces from model (sigma) surfaces." ;
		:platform = "Model" ;
data:

 level = 1000, 925, 850, 700, 600, 500, 400, 300 ;

 lat = 90, 87.5, 85, 82.5, 80, 77.5, 75, 72.5, 70, 67.5, 65, 62.5, 60, 57.5, 
    55, 52.5, 50, 47.5, 45, 42.5, 40, 37.5, 35, 32.5, 30, 27.5, 25, 22.5, 20, 
    17.5, 15, 12.5, 10, 7.5, 5, 2.5, 0, -2.5, -5, -7.5, -10, -12.5, -15, 
    -17.5, -20, -22.5, -25, -27.5, -30, -32.5, -35, -37.5, -40, -42.5, -45, 
    -47.5, -50, -52.5, -55, -57.5, -60, -62.5, -65, -67.5, -70, -72.5, -75, 
    -77.5, -80, -82.5, -85, -87.5, -90 ;

 lon = 0, 2.5, 5, 7.5, 10, 12.5, 15, 17.5, 20, 22.5, 25, 27.5, 30, 32.5, 35, 
    37.5, 40, 42.5, 45, 47.5, 50, 52.5, 55, 57.5, 60, 62.5, 65, 67.5, 70, 
    72.5, 75, 77.5, 80, 82.5, 85, 87.5, 90, 92.5, 95, 97.5, 100, 102.5, 105, 
    107.5, 110, 112.5, 115, 117.5, 120, 122.5, 125, 127.5, 130, 132.5, 135, 
    137.5, 140, 142.5, 145, 147.5, 150, 152.5, 155, 157.5, 160, 162.5, 165, 
    167.5, 170, 172.5, 175, 177.5, 180, 182.5, 185, 187.5, 190, 192.5, 195, 
    197.5, 200, 202.5, 205, 207.5, 210, 212.5, 215, 217.5, 220, 222.5, 225, 
    227.5, 230, 232.5, 235, 237.5, 240, 242.5, 245, 247.5, 250, 252.5, 255, 
    257.5, 260, 262.5, 265, 267.5, 270, 272.5, 275, 277.5, 280, 282.5, 285, 
    287.5, 290, 292.5, 295, 297.5, 300, 302.5, 305, 307.5, 310, 312.5, 315, 
    317.5, 320, 322.5, 325, 327.5, 330, 332.5, 335, 337.5, 340, 342.5, 345, 
    347.5, 350, 352.5, 355, 357.5 ;

 time = 17549208, 17549232, 17549256, 17549280, 17549304, 17549328, 17549352, 
    17549376, 17549400, 17549424, 17549448, 17549472, 17549496, 17549520, 
    17549544, 17549568, 17549592, 17549616, 17549640, 17549664, 17549688, 
    17549712, 17549736, 17549760, 17549784, 17549808, 17549832, 17549856, 
    17549880, 17549904, 17549928, 17549952, 17549976, 17550000, 17550024, 
    17550048, 17550072, 17550096, 17550120, 17550144, 17550168, 17550192, 
    17550216, 17550240, 17550264, 17550288, 17550312, 17550336, 17550360, 
    17550384, 17550408, 17550432, 17550456, 17550480, 17550504, 17550528, 
    17550552, 17550576, 17550600, 17550624, 17550648, 17550672, 17550696, 
    17550720, 17550744, 17550768, 17550792, 17550816, 17550840, 17550864, 
    17550888, 17550912, 17550936, 17550960, 17550984, 17551008, 17551032, 
    17551056, 17551080, 17551104, 17551128, 17551152, 17551176, 17551200, 
    17551224, 17551248, 17551272, 17551296, 17551320, 17551344, 17551368, 
    17551392, 17551416, 17551440, 17551464, 17551488, 17551512, 17551536, 
    17551560, 17551584, 17551608, 17551632, 17551656, 17551680, 17551704, 
    17551728, 17551752, 17551776, 17551800, 17551824, 17551848, 17551872, 
    17551896, 17551920, 17551944, 17551968, 17551992, 17552016, 17552040, 
    17552064, 17552088, 17552112, 17552136, 17552160, 17552184, 17552208, 
    17552232, 17552256, 17552280, 17552304, 17552328, 17552352, 17552376, 
    17552400, 17552424, 17552448, 17552472, 17552496, 17552520, 17552544, 
    17552568, 17552592, 17552616, 17552640, 17552664, 17552688, 17552712, 
    17552736, 17552760, 17552784, 17552808, 17552832, 17552856, 17552880, 
    17552904, 17552928, 17552952, 17552976, 17553000, 17553024, 17553048, 
    17553072, 17553096, 17553120, 17553144, 17553168, 17553192, 17553216, 
    17553240, 17553264, 17553288, 17553312, 17553336, 17553360, 17553384, 
    17553408, 17553432, 17553456, 17553480, 17553504, 17553528, 17553552, 
    17553576, 17553600, 17553624, 17553648, 17553672, 17553696, 17553720, 
    17553744, 17553768, 17553792, 17553816, 17553840, 17553864, 17553888, 
    17553912, 17553936, 17553960, 17553984, 17554008, 17554032, 17554056, 
    17554080, 17554104, 17554128, 17554152, 17554176, 17554200, 17554224, 
    17554248, 17554272, 17554296, 17554320, 17554344, 17554368, 17554392, 
    17554416, 17554440, 17554464, 17554488, 17554512, 17554536, 17554560, 
    17554584, 17554608, 17554632, 17554656, 17554680, 17554704, 17554728, 
    17554752, 17554776, 17554800, 17554824, 17554848, 17554872, 17554896, 
    17554920, 17554944, 17554968, 17554992, 17555016, 17555040, 17555064, 
    17555088, 17555112, 17555136, 17555160, 17555184, 17555208, 17555232, 
    17555256, 17555280, 17555304, 17555328, 17555352, 17555376, 17555400, 
    17555424, 17555448, 17555472, 17555496, 17555520, 17555544, 17555568, 
    17555592, 17555616, 17555640, 17555664, 17555688, 17555712, 17555736, 
    17555760, 17555784, 17555808, 17555832, 17555856, 17555880, 17555904, 
    17555928, 17555952, 17555976, 17556000, 17556024, 17556048, 17556072, 
    17556096, 17556120, 17556144, 17556168, 17556192, 17556216, 17556240, 
    17556264, 17556288, 17556312, 17556336, 17556360, 17556384, 17556408, 
    17556432, 17556456, 17556480, 17556504, 17556528, 17556552, 17556576, 
    17556600, 17556624, 17556648, 17556672, 17556696, 17556720, 17556744, 
    17556768, 17556792, 17556816, 17556840, 17556864, 17556888, 17556912, 
    17556936, 17556960, 17556984, 17557008, 17557032, 17557056, 17557080, 
    17557104, 17557128, 17557152, 17557176, 17557200, 17557224, 17557248, 
    17557272, 17557296, 17557320, 17557344, 17557368, 17557392, 17557416, 
    17557440, 17557464, 17557488, 17557512, 17557536, 17557560, 17557584, 
    17557608, 17557632, 17557656, 17557680, 17557704, 17557728, 17557752, 
    17557776, 17557800, 17557824, 17557848, 17557872, 17557896, 17557920, 
    17557944 ;
}

